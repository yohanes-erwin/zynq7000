// Author: Erwin Ouyang
// Date  : 14 Dec 2018

`timescale 1ns / 1ps

module axi_mm2s_interface
	(
        // ### Clock and reset signals #########################################
        input  wire        aclk,
        input  wire        aresetn,
        // ### AXI4-lite slave signals #########################################
        // *** Write address signals ***
        output wire        s_axi_awready,
        input  wire [31:0] s_axi_awaddr,
        input  wire        s_axi_awvalid,
        // *** Write data signals ***
        output wire        s_axi_wready,
        input  wire [31:0] s_axi_wdata,
        input  wire [3:0]  s_axi_wstrb,
        input  wire        s_axi_wvalid,
        // *** Write response signals ***
        input  wire        s_axi_bready,
        output wire [1:0]  s_axi_bresp,
        output wire        s_axi_bvalid,
        // *** Read address signals ***
        output wire        s_axi_arready,
        input  wire [31:0] s_axi_araddr,
        input  wire        s_axi_arvalid,
        // *** Read data signals ***    
        input  wire        s_axi_rready,
        output wire [31:0] s_axi_rdata,
        output wire [1:0]  s_axi_rresp,
        output wire        s_axi_rvalid,
        // ### AXI4-stream master signals ######################################
        input  wire        m_axis_tready,
        output wire [31:0] m_axis_tdata,
        output wire        m_axis_tvalid,
        output wire        m_axis_tlast,
        // ### User signals ####################################################
        output wire        en,
        output wire [7:0]  mult_const
    );

    // ### Register map ########################################################
    // 0x00: multiplier constant, number of word per frame, enable (active high), and busy
    //       bit 7~0  = CONST[7:0] (R/W)
    //       bit 8~10 = WORD (R/W)
    //       bit 11   = EN (R/W)
    //       bit 12   = BUSY (R)
    // 0x04: data register 0
    //       bit 31~0 = DATA0[31:0] (R/W)
    // 0x08: data register 1
    //       bit 31~0 = DATA1[31:0] (R/W)
    // 0x0c: data register 2
    //       bit 31~0 = DATA2[31:0] (R/W)
    // 0x10: data register 3
    //       bit 31~0 = DATA3[31:0] (R/W)   
	localparam C_ADDR_BITS = 8;
	// *** Address ***
	localparam C_ADDR_CTRL = 8'h00,
			   C_ADDR_DATA0 = 8'h04,
			   C_ADDR_DATA1 = 8'h08,
			   C_ADDR_DATA2 = 8'h0c,
			   C_ADDR_DATA3 = 8'h10;
	// *** AXI write FSM ***
	localparam S_WRIDLE = 2'd0,
			   S_WRDATA = 2'd1,
			   S_WRRESP = 2'd2;
	// *** AXI read FSM ***
	localparam S_RDIDLE = 2'd0,
			   S_RDDATA = 2'd1;
    // *** AXIS FSM ***
    localparam S_IDLE = 2'h0,
               S_WRITE_STREAM = 2'h1;

	// *** AXI write ***
	reg [1:0] wstate_cs, wstate_ns;
	reg [C_ADDR_BITS-1:0] waddr;
	wire [31:0] wmask;
	wire aw_hs, w_hs;
	// *** AXI read ***
	reg [1:0] rstate_cs, rstate_ns;
	wire [C_ADDR_BITS-1:0] raddr;
	reg [31:0] rdata;
	wire ar_hs;
	// *** Control registers ***
    reg [11:0] ctrl_reg;
    wire busy_reg;
    reg [31:0] data_reg [0:3];
    reg start_reg;           
	// *** AXIS ***
    reg [1:0] mm2sstate_cs, mm2sstate_ns;
    reg [1:0] wr_ptr_cv, wr_ptr_nv;
    reg m_axis_tlast_cv, m_axis_tlast_nv;

	// ### AXI write ###########################################################
	assign s_axi_awready = (wstate_cs == S_WRIDLE);
	assign s_axi_wready = (wstate_cs == S_WRDATA);
	assign s_axi_bresp = 2'b00;    // OKAY
	assign s_axi_bvalid = (wstate_cs == S_WRRESP);
	assign wmask = {{8{s_axi_wstrb[3]}}, {8{s_axi_wstrb[2]}}, {8{s_axi_wstrb[1]}}, {8{s_axi_wstrb[0]}}};
	assign aw_hs = s_axi_awvalid & s_axi_awready;
	assign w_hs = s_axi_wvalid & s_axi_wready;

	// *** Write state register ***
	always @(posedge aclk)
	begin
		if (!aresetn)
			wstate_cs <= S_WRIDLE;
		else
			wstate_cs <= wstate_ns;
	end
	
	// *** Write state next ***
	always @(*)
	begin
		case (wstate_cs)
			S_WRIDLE:
				if (s_axi_awvalid)
					wstate_ns = S_WRDATA;
				else
					wstate_ns = S_WRIDLE;
			S_WRDATA:
				if (s_axi_wvalid)
					wstate_ns = S_WRRESP;
				else
					wstate_ns = S_WRDATA;
			S_WRRESP:
				if (s_axi_bready)
					wstate_ns = S_WRIDLE;
				else
					wstate_ns = S_WRRESP;
			default:
				wstate_ns = S_WRIDLE;
		endcase
	end
	
	// *** Write address register ***
	always @(posedge aclk)
	begin
		if (aw_hs)
			waddr <= s_axi_awaddr[C_ADDR_BITS-1:0];
	end   

	// ### AXI read ############################################################
	assign s_axi_arready = (rstate_cs == S_RDIDLE);
	assign s_axi_rdata = rdata;
	assign s_axi_rresp = 2'b00;    // OKAY
	assign s_axi_rvalid = (rstate_cs == S_RDDATA);
	assign ar_hs = s_axi_arvalid & s_axi_arready;
	assign raddr = s_axi_araddr[C_ADDR_BITS-1:0];
	
	// *** Read state register ***
	always @(posedge aclk)
	begin
		if (!aresetn)
			rstate_cs <= S_RDIDLE;
		else
			rstate_cs <= rstate_ns;
	end

	// *** Read state next ***
	always @(*) 
	begin
		case (rstate_cs)
			S_RDIDLE:
				if (s_axi_arvalid)
					rstate_ns = S_RDDATA;
				else
					rstate_ns = S_RDIDLE;
			S_RDDATA:
				if (s_axi_rready)
					rstate_ns = S_RDIDLE;
				else
					rstate_ns = S_RDDATA;
			default:
				rstate_ns = S_RDIDLE;
		endcase
	end
	
	// *** Read data register ***
	always @(posedge aclk)
	begin
	    if (!aresetn)
	        rdata <= 0;
		else if (ar_hs)
			case (raddr)
				C_ADDR_CTRL: 
					rdata <= {busy_reg, ctrl_reg[11:0]};
                C_ADDR_DATA0:
                    rdata <= data_reg[0];
                C_ADDR_DATA1:
                    rdata <= data_reg[1];
                C_ADDR_DATA2:
                    rdata <= data_reg[2];
                C_ADDR_DATA3:
                    rdata <= data_reg[3];   		
			endcase
	end
    
    // ### Control registers ###################################################
   	assign en = ctrl_reg[11]; 
    assign mult_const = ctrl_reg[7:0];
   	
	always @(posedge aclk)
	begin
	    if (!aresetn)
            ctrl_reg[11:0] <= 0;
		else if (w_hs && waddr == C_ADDR_CTRL)
			ctrl_reg[11:0] <= (s_axi_wdata[11:0] & wmask) | (ctrl_reg[11:0] & ~wmask);
	end
	
	always @(posedge aclk)
	begin
	    if (!aresetn)
	    begin
	        start_reg <= 0;
            data_reg[0] <= 0;
            data_reg[1] <= 0;
            data_reg[2] <= 0;
            data_reg[3] <= 0;
        end
		else if (w_hs && waddr == C_ADDR_DATA0)
		begin
		    if (ctrl_reg[10:8] == 1)
                start_reg <= 1;
			data_reg[0][31:0] <= (s_axi_wdata[31:0] & wmask) | (data_reg[0][31:0] & ~wmask);
	    end
		else if (w_hs && waddr == C_ADDR_DATA1)
        begin
            if (ctrl_reg[10:8] == 2)
                start_reg <= 1;
            data_reg[1][31:0] <= (s_axi_wdata[31:0] & wmask) | (data_reg[1][31:0] & ~wmask);
        end
		else if (w_hs && waddr == C_ADDR_DATA2)
        begin
            if (ctrl_reg[10:8] == 3)
                start_reg <= 1;
            data_reg[2][31:0] <= (s_axi_wdata[31:0] & wmask) | (data_reg[2][31:0] & ~wmask);
        end
		else if (w_hs && waddr == C_ADDR_DATA3)
        begin
            if (ctrl_reg[10:8] == 4)
                start_reg <= 1;
            data_reg[3][31:0] <= (s_axi_wdata[31:0] & wmask) | (data_reg[3][31:0] & ~wmask);
        end
	    else
        begin
            start_reg <= 0;
        end
	end

    // ### AXIS ################################################################
    assign busy_reg = (mm2sstate_cs == S_WRITE_STREAM) ? 1 : 0;
    assign m_axis_tdata = data_reg[wr_ptr_cv];
    assign m_axis_tvalid = (mm2sstate_cs == S_WRITE_STREAM) ? 1 : 0;
    assign m_axis_tlast = m_axis_tlast_cv;

    // *** AXIS state register ***
    always @(posedge aclk)
    begin
        if (!aresetn)
        begin
            mm2sstate_cs <= S_IDLE;
            wr_ptr_cv <= 0;
            m_axis_tlast_cv <= 0;
        end
        else
        begin
            mm2sstate_cs <= mm2sstate_ns;
            wr_ptr_cv <= wr_ptr_nv;
            m_axis_tlast_cv <= m_axis_tlast_nv;
        end 
    end

    // *** AXIS state next ***
    always @(*)
    begin
        mm2sstate_ns = mm2sstate_cs;
        wr_ptr_nv = wr_ptr_cv;
        m_axis_tlast_nv = m_axis_tlast_cv;
        case (mm2sstate_cs)
            S_IDLE:
            begin
                if (start_reg)
                begin
                    mm2sstate_ns = S_WRITE_STREAM;
                    if (ctrl_reg[10:8] == 1)
                        m_axis_tlast_nv = 1;    
                end
            end
            S_WRITE_STREAM:
            begin
                if (m_axis_tready)
                begin
                    if (wr_ptr_cv == ctrl_reg[10:8]-1)
                    begin
                        mm2sstate_ns = S_IDLE;
                        wr_ptr_nv = 0;
                        m_axis_tlast_nv = 0;
                    end
                    else
                    begin
                        if (wr_ptr_cv == ctrl_reg[10:8]-2)
                        begin
                            m_axis_tlast_nv = 1;
                        end
                        wr_ptr_nv = wr_ptr_cv + 1;
                    end
                end
            end
        endcase
    end
                         
endmodule
